/***********************************************************************
 * A SystemVerilog testbench for an instruction register.
 * The course labs will convert this to an object-oriented testbench
 * with constrained random test generation, functional coverage, and
 * a scoreboard for self-verification.
 **********************************************************************/

module instr_register_test
  import instr_register_pkg::*;  // user-defined types are defined in instr_register_pkg.sv
  (input  logic          clk,
   output logic          load_en,
   output logic          reset_n,
   output operand_t      operand_a,
   output operand_t      operand_b,
   output opcode_t       opcode,
   output address_t      write_pointer,
   output address_t      read_pointer,
   input  instruction_t  instruction_word
  );

  timeunit 1ns/1ns;

  parameter READ_NR = 9;
  parameter WRITE_NR = 10;

  int seed = 555;

  initial begin
    $display("\n*************************************************************");
    $display(  "***  THIS IS NOW A SELF-CHECKING TESTBENCH. YOU NO        ***");
    $display(  "***  LONGER NEED TO VISUALLY VERIFY THE OUTPUT VALUES     ***");
    $display(  "*** TO MATCH THE INPUT VALUES FOR EACH REGISTER LOCATION  ***");
    $display(  "*************************************************************\n");

    $display("\nReseting the instruction register...");
    write_pointer  = 5'h00;         // initialize write pointer
    read_pointer   = 5'h1F;         // initialize read pointer
    load_en        = 1'b0;          // initialize load control line
    reset_n       <= 1'b0;          // assert reset_n (active low)
    repeat (2) @(posedge clk) ;     // hold in reset for 2 clock cycles
    reset_n        = 1'b1;          // deassert reset_n (active low)

    $display("\nWriting values to register stack...");
    @(posedge clk) load_en = 1'b1;  // enable writing to register
    // repeat (3) begin - 11/03/2024 - GS
    repeat (WRITE_NR) begin
      @(posedge clk) randomize_transaction;
      @(negedge clk) print_transaction;
    end
    @(posedge clk) load_en = 1'b0;  // turn-off writing to register

    // read back and display same three register locations
    $display("\nReading back the same register locations written...");
    // for (int i=0; i<=2; i++) begin - 11/03/2024 - GS
    for (int i=0; i<=READ_NR; i++) begin
      // later labs will replace this loop with iterating through a
      // scoreboard to determine which addresses were written and
      // the expected values to be read back
      @(posedge clk) read_pointer = i;
      @(negedge clk) print_results;
      check_results;
    end

    @(posedge clk) ;
    $display("\n*************************************************************");
    $display(  "***  THIS IS NOW A SELF-CHECKING TESTBENCH. YOU NO        ***");
    $display(  "***  LONGER NEED TO VISUALLY VERIFY THE OUTPUT VALUES     ***");
    $display(  "*** TO MATCH THE INPUT VALUES FOR EACH REGISTER LOCATION  ***");
    $display(  "*************************************************************\n");
    $finish;
  end

  function void randomize_transaction;
    // A later lab will replace this function with SystemVerilog
    // constrained random values
    //
    // The stactic temp variable is required in order to write to fixed
    // addresses of 0, 1 and 2.  This will be replaceed with randomizeed
    // write_pointer values in a later lab
    //
    static int temp = 0;
    operand_a     <= $random(seed)%16;                 // between -15 and 15
    operand_b     <= $unsigned($random)%16;            // between 0 and 15
    opcode        <= opcode_t'($unsigned($random)%8);  // between 0 and 7, cast to opcode_t type
    write_pointer <= temp++;
  endfunction: randomize_transaction

  function void print_transaction;
    $display("Writing to register location %0d: ", write_pointer);
    $display("  opcode = %0d (%s)", opcode, opcode.name);
    $display("  operand_a = %0d",   operand_a);
    $display("  operand_b = %0d\n", operand_b);
  endfunction: print_transaction

  function void print_results;
    $display("Read from register location %0d: ", read_pointer);
    $display("  opcode = %0d (%s)", instruction_word.opc, instruction_word.opc.name);
    $display("  operand_a = %0d",   instruction_word.op_a);
    $display("  operand_b = %0d", instruction_word.op_b);
    $display("  result = %0d\n", instruction_word.res);
  endfunction: print_results

  function void check_results; // din instruction word luam operand A, operand B, op code si calculam iar valorile si le verificam fata de cele din DUT (case)
    automatic longint expected_result = 0; // rezultat intern folosit la calcul, longint e pe 64 de biti, deci pot face comparatie
    if(instruction_word.opc.name == "ZERO")
      expected_result = 0;
    else if(instruction_word.opc.name == "PASSA")
      expected_result = instruction_word.op_a;
    else if(instruction_word.opc.name == "PASSB")
      expected_result = instruction_word.op_b;
    else if(instruction_word.opc.name == "ADD")
      expected_result = instruction_word.op_a + instruction_word.op_b;
    else if(instruction_word.opc.name == "SUB")
      expected_result = instruction_word.op_a - instruction_word.op_b;
    else if(instruction_word.opc.name == "MULT")
      expected_result = instruction_word.op_a * instruction_word.op_b;
    else if(instruction_word.opc.name == "DIV") begin
      if(instruction_word.op_b == 0)
        expected_result = 0;
      else
        expected_result = instruction_word.op_a / instruction_word.op_b;
    end
    else if(instruction_word.opc.name == "MOD")
      expected_result = instruction_word.op_a % instruction_word.op_b;
    
    $display("Read pointer = %0d: ", read_pointer);
    $display("  opcode = %0d (%s)", instruction_word.opc, instruction_word.opc.name);
    $display("  operand_a = %0d",   instruction_word.op_a);
    $display("  operand_b = %0d", instruction_word.op_b);
    $display("  result = %0d", instruction_word.res);
    $display("  expected result = %0d", expected_result);
    
    if(expected_result == instruction_word.res)
      $display("OK: Expected result and the actual result are identical!\n");
    else
      $display("ERROR: Expected result and the actual result differ!\n");
  endfunction: check_results

endmodule: instr_register_test
